`timescale 1 ns / 1 ps

module AESL_deadlock_kernel_monitor_top ( 
    input wire kernel_monitor_clock,
    input wire kernel_monitor_reset
);
wire [1:0] axis_block_sigs;
wire [17:0] inst_idle_sigs;
wire [13:0] inst_block_sigs;
wire kernel_block;

assign axis_block_sigs[0] = ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.input_layer_TDATA_blk_n;
assign axis_block_sigs[1] = ~AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.grp_softmax_stable_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_s_fu_26.layer21_out_TDATA_blk_n;

assign inst_idle_sigs[0] = AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.ap_idle;
assign inst_block_sigs[0] = (AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.ap_done & ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.ap_continue) | ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.layer2_out_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_22_14_5_3_0_6u_config2_s_fu_116.layer2_out_blk_n;
assign inst_idle_sigs[1] = AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_6u_hard_tanh_config4_U0.ap_idle;
assign inst_block_sigs[1] = (AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_6u_hard_tanh_config4_U0.ap_done & ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_6u_hard_tanh_config4_U0.ap_continue) | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_6u_hard_tanh_config4_U0.layer2_out_blk_n | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_6u_hard_tanh_config4_U0.layer4_out_blk_n;
assign inst_idle_sigs[2] = AESL_inst_myproject.pooling2d_cl_array_ap_fixed_6u_array_ap_fixed_8_1_4_0_0_6u_config5_U0.ap_idle;
assign inst_block_sigs[2] = (AESL_inst_myproject.pooling2d_cl_array_ap_fixed_6u_array_ap_fixed_8_1_4_0_0_6u_config5_U0.ap_done & ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_6u_array_ap_fixed_8_1_4_0_0_6u_config5_U0.ap_continue) | ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_6u_array_ap_fixed_8_1_4_0_0_6u_config5_U0.layer4_out_blk_n | ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_6u_array_ap_fixed_8_1_4_0_0_6u_config5_U0.layer5_out_blk_n;
assign inst_idle_sigs[3] = AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.ap_idle;
assign inst_block_sigs[3] = (AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.ap_done & ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.ap_continue) | ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.layer5_out_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.layer6_out_blk_n | ~AESL_inst_myproject.conv_2d_cl_array_ap_fixed_6u_array_ap_fixed_25_14_5_3_0_16u_config6_U0.grp_compute_output_buffer_2d_array_array_ap_fixed_25_14_5_3_0_16u_config6_s_fu_424.layer6_out_blk_n;
assign inst_idle_sigs[4] = AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config8_U0.ap_idle;
assign inst_block_sigs[4] = (AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config8_U0.ap_done & ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config8_U0.ap_continue) | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config8_U0.layer6_out_blk_n | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config8_U0.layer8_out_blk_n;
assign inst_idle_sigs[5] = AESL_inst_myproject.pooling2d_cl_array_ap_fixed_16u_array_ap_fixed_8_1_4_0_0_16u_config9_U0.ap_idle;
assign inst_block_sigs[5] = (AESL_inst_myproject.pooling2d_cl_array_ap_fixed_16u_array_ap_fixed_8_1_4_0_0_16u_config9_U0.ap_done & ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_16u_array_ap_fixed_8_1_4_0_0_16u_config9_U0.ap_continue) | ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_16u_array_ap_fixed_8_1_4_0_0_16u_config9_U0.layer8_out_blk_n | ~AESL_inst_myproject.pooling2d_cl_array_ap_fixed_16u_array_ap_fixed_8_1_4_0_0_16u_config9_U0.layer9_out_blk_n;
assign inst_idle_sigs[6] = AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_25_14_5_3_0_16u_config11_U0.ap_idle;
assign inst_block_sigs[6] = (AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_25_14_5_3_0_16u_config11_U0.ap_done & ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_25_14_5_3_0_16u_config11_U0.ap_continue) | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_25_14_5_3_0_16u_config11_U0.grp_dense_array_array_ap_fixed_25_14_5_3_0_16u_config11_Pipeline_DataPrepare_fu_1057.layer9_out_blk_n | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_25_14_5_3_0_16u_config11_U0.layer11_out_blk_n;
assign inst_idle_sigs[7] = AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_34_19_5_3_0_16u_config13_U0.ap_idle;
assign inst_block_sigs[7] = (AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_34_19_5_3_0_16u_config13_U0.ap_done & ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_34_19_5_3_0_16u_config13_U0.ap_continue) | ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_34_19_5_3_0_16u_config13_U0.layer11_out_blk_n | ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_34_19_5_3_0_16u_config13_U0.layer13_out_blk_n;
assign inst_idle_sigs[8] = AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config14_U0.ap_idle;
assign inst_block_sigs[8] = (AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config14_U0.ap_done & ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config14_U0.ap_continue) | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config14_U0.layer13_out_blk_n | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config14_U0.layer14_out_blk_n;
assign inst_idle_sigs[9] = AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_16u_config15_U0.ap_idle;
assign inst_block_sigs[9] = (AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_16u_config15_U0.ap_done & ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_16u_config15_U0.ap_continue) | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_16u_config15_U0.layer14_out_blk_n | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_16u_config15_U0.layer15_out_blk_n;
assign inst_idle_sigs[10] = AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_30_15_5_3_0_16u_config17_U0.ap_idle;
assign inst_block_sigs[10] = (AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_30_15_5_3_0_16u_config17_U0.ap_done & ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_30_15_5_3_0_16u_config17_U0.ap_continue) | ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_30_15_5_3_0_16u_config17_U0.layer15_out_blk_n | ~AESL_inst_myproject.normalize_array_ap_fixed_16u_array_ap_fixed_30_15_5_3_0_16u_config17_U0.layer17_out_blk_n;
assign inst_idle_sigs[11] = AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config18_U0.ap_idle;
assign inst_block_sigs[11] = (AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config18_U0.ap_done & ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config18_U0.ap_continue) | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config18_U0.layer17_out_blk_n | ~AESL_inst_myproject.hard_tanh_array_array_ap_fixed_8_1_4_0_0_16u_hard_tanh_config18_U0.layer18_out_blk_n;
assign inst_idle_sigs[12] = AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_10u_config19_U0.ap_idle;
assign inst_block_sigs[12] = (AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_10u_config19_U0.ap_done & ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_10u_config19_U0.ap_continue) | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_10u_config19_U0.layer18_out_blk_n | ~AESL_inst_myproject.dense_array_ap_fixed_16u_array_ap_fixed_21_10_5_3_0_10u_config19_U0.layer19_out_blk_n;
assign inst_idle_sigs[13] = AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.ap_idle;
assign inst_block_sigs[13] = (AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.ap_done & ~AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.ap_continue) | ~AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.grp_softmax_stable_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_s_fu_26.layer19_out_blk_n;

assign inst_idle_sigs[14] = 1'b0;
assign inst_idle_sigs[15] = AESL_inst_myproject.conv_2d_cl_array_ap_fixed_1u_array_ap_fixed_22_14_5_3_0_6u_config2_U0.ap_idle;
assign inst_idle_sigs[16] = AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.ap_idle;
assign inst_idle_sigs[17] = AESL_inst_myproject.softmax_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_U0.grp_softmax_stable_array_array_ap_fixed_8_4_5_3_0_10u_softmax_config21_s_fu_26.ap_idle;

AESL_deadlock_idx0_monitor AESL_deadlock_idx0_monitor_U (
    .clock(kernel_monitor_clock),
    .reset(kernel_monitor_reset),
    .axis_block_sigs(axis_block_sigs),
    .inst_idle_sigs(inst_idle_sigs),
    .inst_block_sigs(inst_block_sigs),
    .block(kernel_block)
);


initial begin : trigger_axis_deadlock
reg block_delay;
    block_delay = 0;
    while(1) begin
        @(posedge kernel_monitor_clock);
    if (kernel_block == 1'b1 && block_delay == 1'b0)
        block_delay = kernel_block;
    end
end

endmodule
